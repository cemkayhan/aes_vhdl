library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_lib.BYTE;

entity multiply_d is
	port (i : in BYTE;
			o : out BYTE
			);
			
end multiply_d;

architecture Behavioral of multiply_d is

begin
	with i select o <=
		x"00" when x"00",
		x"0D" when x"01",
		x"1A" when x"02",
		x"17" when x"03",
		x"34" when x"04",
		x"39" when x"05",
		x"2E" when x"06",
		x"23" when x"07",
		x"68" when x"08",
		x"65" when x"09",
		x"72" when x"0A",
		x"7F" when x"0B",
		x"5C" when x"0C",
		x"51" when x"0D",
		x"46" when x"0E",
		x"4B" when x"0F",
		x"D0" when x"10",
		x"DD" when x"11",
		x"CA" when x"12",
		x"C7" when x"13",
		x"E4" when x"14",
		x"E9" when x"15",
		x"FE" when x"16",
		x"F3" when x"17",
		x"B8" when x"18",
		x"B5" when x"19",
		x"A2" when x"1A",
		x"AF" when x"1B",
		x"8C" when x"1C",
		x"81" when x"1D",
		x"96" when x"1E",
		x"9B" when x"1F",
		x"BB" when x"20",
		x"B6" when x"21",
		x"A1" when x"22",
		x"AC" when x"23",
		x"8F" when x"24",
		x"82" when x"25",
		x"95" when x"26",
		x"98" when x"27",
		x"D3" when x"28",
		x"DE" when x"29",
		x"C9" when x"2A",
		x"C4" when x"2B",
		x"E7" when x"2C",
		x"EA" when x"2D",
		x"FD" when x"2E",
		x"F0" when x"2F",
		x"6B" when x"30",
		x"66" when x"31",
		x"71" when x"32",
		x"7C" when x"33",
		x"5F" when x"34",
		x"52" when x"35",
		x"45" when x"36",
		x"48" when x"37",
		x"03" when x"38",
		x"0E" when x"39",
		x"19" when x"3A",
		x"14" when x"3B",
		x"37" when x"3C",
		x"3A" when x"3D",
		x"2D" when x"3E",
		x"20" when x"3F",
		x"6D" when x"40",
		x"60" when x"41",
		x"77" when x"42",
		x"7A" when x"43",
		x"59" when x"44",
		x"54" when x"45",
		x"43" when x"46",
		x"4E" when x"47",
		x"05" when x"48",
		x"08" when x"49",
		x"1F" when x"4A",
		x"12" when x"4B",
		x"31" when x"4C",
		x"3C" when x"4D",
		x"2B" when x"4E",
		x"26" when x"4F",
		x"BD" when x"50",
		x"B0" when x"51",
		x"A7" when x"52",
		x"AA" when x"53",
		x"89" when x"54",
		x"84" when x"55",
		x"93" when x"56",
		x"9E" when x"57",
		x"D5" when x"58",
		x"D8" when x"59",
		x"CF" when x"5A",
		x"C2" when x"5B",
		x"E1" when x"5C",
		x"EC" when x"5D",
		x"FB" when x"5E",
		x"F6" when x"5F",
		x"D6" when x"60",
		x"DB" when x"61",
		x"CC" when x"62",
		x"C1" when x"63",
		x"E2" when x"64",
		x"EF" when x"65",
		x"F8" when x"66",
		x"F5" when x"67",
		x"BE" when x"68",
		x"B3" when x"69",
		x"A4" when x"6A",
		x"A9" when x"6B",
		x"8A" when x"6C",
		x"87" when x"6D",
		x"90" when x"6E",
		x"9D" when x"6F",
		x"06" when x"70",
		x"0B" when x"71",
		x"1C" when x"72",
		x"11" when x"73",
		x"32" when x"74",
		x"3F" when x"75",
		x"28" when x"76",
		x"25" when x"77",
		x"6E" when x"78",
		x"63" when x"79",
		x"74" when x"7A",
		x"79" when x"7B",
		x"5A" when x"7C",
		x"57" when x"7D",
		x"40" when x"7E",
		x"4D" when x"7F",
		x"DA" when x"80",
		x"D7" when x"81",
		x"C0" when x"82",
		x"CD" when x"83",
		x"EE" when x"84",
		x"E3" when x"85",
		x"F4" when x"86",
		x"F9" when x"87",
		x"B2" when x"88",
		x"BF" when x"89",
		x"A8" when x"8A",
		x"A5" when x"8B",
		x"86" when x"8C",
		x"8B" when x"8D",
		x"9C" when x"8E",
		x"91" when x"8F",
		x"0A" when x"90",
		x"07" when x"91",
		x"10" when x"92",
		x"1D" when x"93",
		x"3E" when x"94",
		x"33" when x"95",
		x"24" when x"96",
		x"29" when x"97",
		x"62" when x"98",
		x"6F" when x"99",
		x"78" when x"9A",
		x"75" when x"9B",
		x"56" when x"9C",
		x"5B" when x"9D",
		x"4C" when x"9E",
		x"41" when x"9F",
		x"61" when x"A0",
		x"6C" when x"A1",
		x"7B" when x"A2",
		x"76" when x"A3",
		x"55" when x"A4",
		x"58" when x"A5",
		x"4F" when x"A6",
		x"42" when x"A7",
		x"09" when x"A8",
		x"04" when x"A9",
		x"13" when x"AA",
		x"1E" when x"AB",
		x"3D" when x"AC",
		x"30" when x"AD",
		x"27" when x"AE",
		x"2A" when x"AF",
		x"B1" when x"B0",
		x"BC" when x"B1",
		x"AB" when x"B2",
		x"A6" when x"B3",
		x"85" when x"B4",
		x"88" when x"B5",
		x"9F" when x"B6",
		x"92" when x"B7",
		x"D9" when x"B8",
		x"D4" when x"B9",
		x"C3" when x"BA",
		x"CE" when x"BB",
		x"ED" when x"BC",
		x"E0" when x"BD",
		x"F7" when x"BE",
		x"FA" when x"BF",
		x"B7" when x"C0",
		x"BA" when x"C1",
		x"AD" when x"C2",
		x"A0" when x"C3",
		x"83" when x"C4",
		x"8E" when x"C5",
		x"99" when x"C6",
		x"94" when x"C7",
		x"DF" when x"C8",
		x"D2" when x"C9",
		x"C5" when x"CA",
		x"C8" when x"CB",
		x"EB" when x"CC",
		x"E6" when x"CD",
		x"F1" when x"CE",
		x"FC" when x"CF",
		x"67" when x"D0",
		x"6A" when x"D1",
		x"7D" when x"D2",
		x"70" when x"D3",
		x"53" when x"D4",
		x"5E" when x"D5",
		x"49" when x"D6",
		x"44" when x"D7",
		x"0F" when x"D8",
		x"02" when x"D9",
		x"15" when x"DA",
		x"18" when x"DB",
		x"3B" when x"DC",
		x"36" when x"DD",
		x"21" when x"DE",
		x"2C" when x"DF",
		x"0C" when x"E0",
		x"01" when x"E1",
		x"16" when x"E2",
		x"1B" when x"E3",
		x"38" when x"E4",
		x"35" when x"E5",
		x"22" when x"E6",
		x"2F" when x"E7",
		x"64" when x"E8",
		x"69" when x"E9",
		x"7E" when x"EA",
		x"73" when x"EB",
		x"50" when x"EC",
		x"5D" when x"ED",
		x"4A" when x"EE",
		x"47" when x"EF",
		x"DC" when x"F0",
		x"D1" when x"F1",
		x"C6" when x"F2",
		x"CB" when x"F3",
		x"E8" when x"F4",
		x"E5" when x"F5",
		x"F2" when x"F6",
		x"FF" when x"F7",
		x"B4" when x"F8",
		x"B9" when x"F9",
		x"AE" when x"FA",
		x"A3" when x"FB",
		x"80" when x"FC",
		x"8D" when x"FD",
		x"9A" when x"FE",
		x"97" when x"FF",
		x"00" when others;

end Behavioral;

