library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_lib.BYTE;

entity multiply_9 is
	port (i : in BYTE;
			o : out BYTE
			);
			
end multiply_9;

architecture Behavioral of multiply_9 is

begin
	with i select o <=
		x"00" when x"00",
		x"09" when x"01",
		x"12" when x"02",
		x"1B" when x"03",
		x"24" when x"04",
		x"2D" when x"05",
		x"36" when x"06",
		x"3F" when x"07",
		x"48" when x"08",
		x"41" when x"09",
		x"5A" when x"0A",
		x"53" when x"0B",
		x"6C" when x"0C",
		x"65" when x"0D",
		x"7E" when x"0E",
		x"77" when x"0F",
		x"90" when x"10",
		x"99" when x"11",
		x"82" when x"12",
		x"8B" when x"13",
		x"B4" when x"14",
		x"BD" when x"15",
		x"A6" when x"16",
		x"AF" when x"17",
		x"D8" when x"18",
		x"D1" when x"19",
		x"CA" when x"1A",
		x"C3" when x"1B",
		x"FC" when x"1C",
		x"F5" when x"1D",
		x"EE" when x"1E",
		x"E7" when x"1F",
		x"3B" when x"20",
		x"32" when x"21",
		x"29" when x"22",
		x"20" when x"23",
		x"1F" when x"24",
		x"16" when x"25",
		x"0D" when x"26",
		x"04" when x"27",
		x"73" when x"28",
		x"7A" when x"29",
		x"61" when x"2A",
		x"68" when x"2B",
		x"57" when x"2C",
		x"5E" when x"2D",
		x"45" when x"2E",
		x"4C" when x"2F",
		x"AB" when x"30",
		x"A2" when x"31",
		x"B9" when x"32",
		x"B0" when x"33",
		x"8F" when x"34",
		x"86" when x"35",
		x"9D" when x"36",
		x"94" when x"37",
		x"E3" when x"38",
		x"EA" when x"39",
		x"F1" when x"3A",
		x"F8" when x"3B",
		x"C7" when x"3C",
		x"CE" when x"3D",
		x"D5" when x"3E",
		x"DC" when x"3F",
		x"76" when x"40",
		x"7F" when x"41",
		x"64" when x"42",
		x"6D" when x"43",
		x"52" when x"44",
		x"5B" when x"45",
		x"40" when x"46",
		x"49" when x"47",
		x"3E" when x"48",
		x"37" when x"49",
		x"2C" when x"4A",
		x"25" when x"4B",
		x"1A" when x"4C",
		x"13" when x"4D",
		x"08" when x"4E",
		x"01" when x"4F",
		x"E6" when x"50",
		x"EF" when x"51",
		x"F4" when x"52",
		x"FD" when x"53",
		x"C2" when x"54",
		x"CB" when x"55",
		x"D0" when x"56",
		x"D9" when x"57",
		x"AE" when x"58",
		x"A7" when x"59",
		x"BC" when x"5A",
		x"B5" when x"5B",
		x"8A" when x"5C",
		x"83" when x"5D",
		x"98" when x"5E",
		x"91" when x"5F",
		x"4D" when x"60",
		x"44" when x"61",
		x"5F" when x"62",
		x"56" when x"63",
		x"69" when x"64",
		x"60" when x"65",
		x"7B" when x"66",
		x"72" when x"67",
		x"05" when x"68",
		x"0C" when x"69",
		x"17" when x"6A",
		x"1E" when x"6B",
		x"21" when x"6C",
		x"28" when x"6D",
		x"33" when x"6E",
		x"3A" when x"6F",
		x"DD" when x"70",
		x"D4" when x"71",
		x"CF" when x"72",
		x"C6" when x"73",
		x"F9" when x"74",
		x"F0" when x"75",
		x"EB" when x"76",
		x"E2" when x"77",
		x"95" when x"78",
		x"9C" when x"79",
		x"87" when x"7A",
		x"8E" when x"7B",
		x"B1" when x"7C",
		x"B8" when x"7D",
		x"A3" when x"7E",
		x"AA" when x"7F",
		x"EC" when x"80",
		x"E5" when x"81",
		x"FE" when x"82",
		x"F7" when x"83",
		x"C8" when x"84",
		x"C1" when x"85",
		x"DA" when x"86",
		x"D3" when x"87",
		x"A4" when x"88",
		x"AD" when x"89",
		x"B6" when x"8A",
		x"BF" when x"8B",
		x"80" when x"8C",
		x"89" when x"8D",
		x"92" when x"8E",
		x"9B" when x"8F",
		x"7C" when x"90",
		x"75" when x"91",
		x"6E" when x"92",
		x"67" when x"93",
		x"58" when x"94",
		x"51" when x"95",
		x"4A" when x"96",
		x"43" when x"97",
		x"34" when x"98",
		x"3D" when x"99",
		x"26" when x"9A",
		x"2F" when x"9B",
		x"10" when x"9C",
		x"19" when x"9D",
		x"02" when x"9E",
		x"0B" when x"9F",
		x"D7" when x"A0",
		x"DE" when x"A1",
		x"C5" when x"A2",
		x"CC" when x"A3",
		x"F3" when x"A4",
		x"FA" when x"A5",
		x"E1" when x"A6",
		x"E8" when x"A7",
		x"9F" when x"A8",
		x"96" when x"A9",
		x"8D" when x"AA",
		x"84" when x"AB",
		x"BB" when x"AC",
		x"B2" when x"AD",
		x"A9" when x"AE",
		x"A0" when x"AF",
		x"47" when x"B0",
		x"4E" when x"B1",
		x"55" when x"B2",
		x"5C" when x"B3",
		x"63" when x"B4",
		x"6A" when x"B5",
		x"71" when x"B6",
		x"78" when x"B7",
		x"0F" when x"B8",
		x"06" when x"B9",
		x"1D" when x"BA",
		x"14" when x"BB",
		x"2B" when x"BC",
		x"22" when x"BD",
		x"39" when x"BE",
		x"30" when x"BF",
		x"9A" when x"C0",
		x"93" when x"C1",
		x"88" when x"C2",
		x"81" when x"C3",
		x"BE" when x"C4",
		x"B7" when x"C5",
		x"AC" when x"C6",
		x"A5" when x"C7",
		x"D2" when x"C8",
		x"DB" when x"C9",
		x"C0" when x"CA",
		x"C9" when x"CB",
		x"F6" when x"CC",
		x"FF" when x"CD",
		x"E4" when x"CE",
		x"ED" when x"CF",
		x"0A" when x"D0",
		x"03" when x"D1",
		x"18" when x"D2",
		x"11" when x"D3",
		x"2E" when x"D4",
		x"27" when x"D5",
		x"3C" when x"D6",
		x"35" when x"D7",
		x"42" when x"D8",
		x"4B" when x"D9",
		x"50" when x"DA",
		x"59" when x"DB",
		x"66" when x"DC",
		x"6F" when x"DD",
		x"74" when x"DE",
		x"7D" when x"DF",
		x"A1" when x"E0",
		x"A8" when x"E1",
		x"B3" when x"E2",
		x"BA" when x"E3",
		x"85" when x"E4",
		x"8C" when x"E5",
		x"97" when x"E6",
		x"9E" when x"E7",
		x"E9" when x"E8",
		x"E0" when x"E9",
		x"FB" when x"EA",
		x"F2" when x"EB",
		x"CD" when x"EC",
		x"C4" when x"ED",
		x"DF" when x"EE",
		x"D6" when x"EF",
		x"31" when x"F0",
		x"38" when x"F1",
		x"23" when x"F2",
		x"2A" when x"F3",
		x"15" when x"F4",
		x"1C" when x"F5",
		x"07" when x"F6",
		x"0E" when x"F7",
		x"79" when x"F8",
		x"70" when x"F9",
		x"6B" when x"FA",
		x"62" when x"FB",
		x"5D" when x"FC",
		x"54" when x"FD",
		x"4F" when x"FE",
		x"46" when x"FF",
		x"00" when others;  

end Behavioral;

