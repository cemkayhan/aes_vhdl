library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiply_e is
	port (i : in std_logic_vector (7 downto 0);
			o : out std_logic_vector (7 downto 0)
			);
			
end multiply_e;

architecture Behavioral of multiply_e is
	
begin
	with i select o <=
		x"00" when x"00",
		x"0E" when x"01",
		x"1C" when x"02",
		x"12" when x"03",
		x"38" when x"04",
		x"36" when x"05",
		x"24" when x"06",
		x"2A" when x"07",
		x"70" when x"08",
		x"7E" when x"09",
		x"6C" when x"0A",
		x"62" when x"0B",
		x"48" when x"0C",
		x"46" when x"0D",
		x"54" when x"0E",
		x"5A" when x"0F",
		x"E0" when x"10",
		x"EE" when x"11",
		x"FC" when x"12",
		x"F2" when x"13",
		x"D8" when x"14",
		x"D6" when x"15",
		x"C4" when x"16",
		x"CA" when x"17",
		x"90" when x"18",
		x"9E" when x"19",
		x"8C" when x"1A",
		x"82" when x"1B",
		x"A8" when x"1C",
		x"A6" when x"1D",
		x"B4" when x"1E",
		x"BA" when x"1F",
		x"DB" when x"20",
		x"D5" when x"21",
		x"C7" when x"22",
		x"C9" when x"23",
		x"E3" when x"24",
		x"ED" when x"25",
		x"FF" when x"26",
		x"F1" when x"27",
		x"AB" when x"28",
		x"A5" when x"29",
		x"B7" when x"2A",
		x"B9" when x"2B",
		x"93" when x"2C",
		x"9D" when x"2D",
		x"8F" when x"2E",
		x"81" when x"2F",
		x"3B" when x"30",
		x"35" when x"31",
		x"27" when x"32",
		x"29" when x"33",
		x"03" when x"34",
		x"0D" when x"35",
		x"1F" when x"36",
		x"11" when x"37",
		x"4B" when x"38",
		x"45" when x"39",
		x"57" when x"3A",
		x"59" when x"3B",
		x"73" when x"3C",
		x"7D" when x"3D",
		x"6F" when x"3E",
		x"61" when x"3F",
		x"AD" when x"40",
		x"A3" when x"41",
		x"B1" when x"42",
		x"BF" when x"43",
		x"95" when x"44",
		x"9B" when x"45",
		x"89" when x"46",
		x"87" when x"47",
		x"DD" when x"48",
		x"D3" when x"49",
		x"C1" when x"4A",
		x"CF" when x"4B",
		x"E5" when x"4C",
		x"EB" when x"4D",
		x"F9" when x"4E",
		x"F7" when x"4F",
		x"4D" when x"50",
		x"43" when x"51",
		x"51" when x"52",
		x"5F" when x"53",
		x"75" when x"54",
		x"7B" when x"55",
		x"69" when x"56",
		x"67" when x"57",
		x"3D" when x"58",
		x"33" when x"59",
		x"21" when x"5A",
		x"2F" when x"5B",
		x"05" when x"5C",
		x"0B" when x"5D",
		x"19" when x"5E",
		x"17" when x"5F",
		x"76" when x"60",
		x"78" when x"61",
		x"6A" when x"62",
		x"64" when x"63",
		x"4E" when x"64",
		x"40" when x"65",
		x"52" when x"66",
		x"5C" when x"67",
		x"06" when x"68",
		x"08" when x"69",
		x"1A" when x"6A",
		x"14" when x"6B",
		x"3E" when x"6C",
		x"30" when x"6D",
		x"22" when x"6E",
		x"2C" when x"6F",
		x"96" when x"70",
		x"98" when x"71",
		x"8A" when x"72",
		x"84" when x"73",
		x"AE" when x"74",
		x"A0" when x"75",
		x"B2" when x"76",
		x"BC" when x"77",
		x"E6" when x"78",
		x"E8" when x"79",
		x"FA" when x"7A",
		x"F4" when x"7B",
		x"DE" when x"7C",
		x"D0" when x"7D",
		x"C2" when x"7E",
		x"CC" when x"7F",
		x"41" when x"80",
		x"4F" when x"81",
		x"5D" when x"82",
		x"53" when x"83",
		x"79" when x"84",
		x"77" when x"85",
		x"65" when x"86",
		x"6B" when x"87",
		x"31" when x"88",
		x"3F" when x"89",
		x"2D" when x"8A",
		x"23" when x"8B",
		x"09" when x"8C",
		x"07" when x"8D",
		x"15" when x"8E",
		x"1B" when x"8F",
		x"A1" when x"90",
		x"AF" when x"91",
		x"BD" when x"92",
		x"B3" when x"93",
		x"99" when x"94",
		x"97" when x"95",
		x"85" when x"96",
		x"8B" when x"97",
		x"D1" when x"98",
		x"DF" when x"99",
		x"CD" when x"9A",
		x"C3" when x"9B",
		x"E9" when x"9C",
		x"E7" when x"9D",
		x"F5" when x"9E",
		x"FB" when x"9F",
		x"9A" when x"A0",
		x"94" when x"A1",
		x"86" when x"A2",
		x"88" when x"A3",
		x"A2" when x"A4",
		x"AC" when x"A5",
		x"BE" when x"A6",
		x"B0" when x"A7",
		x"EA" when x"A8",
		x"E4" when x"A9",
		x"F6" when x"AA",
		x"F8" when x"AB",
		x"D2" when x"AC",
		x"DC" when x"AD",
		x"CE" when x"AE",
		x"C0" when x"AF",
		x"7A" when x"B0",
		x"74" when x"B1",
		x"66" when x"B2",
		x"68" when x"B3",
		x"42" when x"B4",
		x"4C" when x"B5",
		x"5E" when x"B6",
		x"50" when x"B7",
		x"0A" when x"B8",
		x"04" when x"B9",
		x"16" when x"BA",
		x"18" when x"BB",
		x"32" when x"BC",
		x"3C" when x"BD",
		x"2E" when x"BE",
		x"20" when x"BF",
		x"EC" when x"C0",
		x"E2" when x"C1",
		x"F0" when x"C2",
		x"FE" when x"C3",
		x"D4" when x"C4",
		x"DA" when x"C5",
		x"C8" when x"C6",
		x"C6" when x"C7",
		x"9C" when x"C8",
		x"92" when x"C9",
		x"80" when x"CA",
		x"8E" when x"CB",
		x"A4" when x"CC",
		x"AA" when x"CD",
		x"B8" when x"CE",
		x"B6" when x"CF",
		x"0C" when x"D0",
		x"02" when x"D1",
		x"10" when x"D2",
		x"1E" when x"D3",
		x"34" when x"D4",
		x"3A" when x"D5",
		x"28" when x"D6",
		x"26" when x"D7",
		x"7C" when x"D8",
		x"72" when x"D9",
		x"60" when x"DA",
		x"6E" when x"DB",
		x"44" when x"DC",
		x"4A" when x"DD",
		x"58" when x"DE",
		x"56" when x"DF",
		x"37" when x"E0",
		x"39" when x"E1",
		x"2B" when x"E2",
		x"25" when x"E3",
		x"0F" when x"E4",
		x"01" when x"E5",
		x"13" when x"E6",
		x"1D" when x"E7",
		x"47" when x"E8",
		x"49" when x"E9",
		x"5B" when x"EA",
		x"55" when x"EB",
		x"7F" when x"EC",
		x"71" when x"ED",
		x"63" when x"EE",
		x"6D" when x"EF",
		x"D7" when x"F0",
		x"D9" when x"F1",
		x"CB" when x"F2",
		x"C5" when x"F3",
		x"EF" when x"F4",
		x"E1" when x"F5",
		x"F3" when x"F6",
		x"FD" when x"F7",
		x"A7" when x"F8",
		x"A9" when x"F9",
		x"BB" when x"FA",
		x"B5" when x"FB",
		x"9F" when x"FC",
		x"91" when x"FD",
		x"83" when x"FE",
		x"8D" when x"FF",
		x"00" when others;  

end Behavioral;

