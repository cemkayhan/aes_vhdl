library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.aes_lib.BYTE;

entity multiply_2 is
	port (i : in BYTE;
			o : out BYTE
			);
			
end multiply_2;

architecture Behavioral of multiply_2 is

begin
	with i select o <=
		x"00" when x"00",
		x"02" when x"01",
		x"04" when x"02",
		x"06" when x"03",
		x"08" when x"04",
		x"0A" when x"05",
		x"0C" when x"06",
		x"0E" when x"07",
		x"10" when x"08",
		x"12" when x"09",
		x"14" when x"0A",
		x"16" when x"0B",
		x"18" when x"0C",
		x"1A" when x"0D",
		x"1C" when x"0E",
		x"1E" when x"0F",
		x"20" when x"10",
		x"22" when x"11",
		x"24" when x"12",
		x"26" when x"13",
		x"28" when x"14",
		x"2A" when x"15",
		x"2C" when x"16",
		x"2E" when x"17",
		x"30" when x"18",
		x"32" when x"19",
		x"34" when x"1A",
		x"36" when x"1B",
		x"38" when x"1C",
		x"3A" when x"1D",
		x"3C" when x"1E",
		x"3E" when x"1F",
		x"40" when x"20",
		x"42" when x"21",
		x"44" when x"22",
		x"46" when x"23",
		x"48" when x"24",
		x"4A" when x"25",
		x"4C" when x"26",
		x"4E" when x"27",
		x"50" when x"28",
		x"52" when x"29",
		x"54" when x"2A",
		x"56" when x"2B",
		x"58" when x"2C",
		x"5A" when x"2D",
		x"5C" when x"2E",
		x"5E" when x"2F",
		x"60" when x"30",
		x"62" when x"31",
		x"64" when x"32",
		x"66" when x"33",
		x"68" when x"34",
		x"6A" when x"35",
		x"6C" when x"36",
		x"6E" when x"37",
		x"70" when x"38",
		x"72" when x"39",
		x"74" when x"3A",
		x"76" when x"3B",
		x"78" when x"3C",
		x"7A" when x"3D",
		x"7C" when x"3E",
		x"7E" when x"3F",
		x"80" when x"40",
		x"82" when x"41",
		x"84" when x"42",
		x"86" when x"43",
		x"88" when x"44",
		x"8A" when x"45",
		x"8C" when x"46",
		x"8E" when x"47",
		x"90" when x"48",
		x"92" when x"49",
		x"94" when x"4A",
		x"96" when x"4B",
		x"98" when x"4C",
		x"9A" when x"4D",
		x"9C" when x"4E",
		x"9E" when x"4F",
		x"A0" when x"50",
		x"A2" when x"51",
		x"A4" when x"52",
		x"A6" when x"53",
		x"A8" when x"54",
		x"AA" when x"55",
		x"AC" when x"56",
		x"AE" when x"57",
		x"B0" when x"58",
		x"B2" when x"59",
		x"B4" when x"5A",
		x"B6" when x"5B",
		x"B8" when x"5C",
		x"BA" when x"5D",
		x"BC" when x"5E",
		x"BE" when x"5F",
		x"C0" when x"60",
		x"C2" when x"61",
		x"C4" when x"62",
		x"C6" when x"63",
		x"C8" when x"64",
		x"CA" when x"65",
		x"CC" when x"66",
		x"CE" when x"67",
		x"D0" when x"68",
		x"D2" when x"69",
		x"D4" when x"6A",
		x"D6" when x"6B",
		x"D8" when x"6C",
		x"DA" when x"6D",
		x"DC" when x"6E",
		x"DE" when x"6F",
		x"E0" when x"70",
		x"E2" when x"71",
		x"E4" when x"72",
		x"E6" when x"73",
		x"E8" when x"74",
		x"EA" when x"75",
		x"EC" when x"76",
		x"EE" when x"77",
		x"F0" when x"78",
		x"F2" when x"79",
		x"F4" when x"7A",
		x"F6" when x"7B",
		x"F8" when x"7C",
		x"FA" when x"7D",
		x"FC" when x"7E",
		x"FE" when x"7F",
		x"1B" when x"80",
		x"19" when x"81",
		x"1F" when x"82",
		x"1D" when x"83",
		x"13" when x"84",
		x"11" when x"85",
		x"17" when x"86",
		x"15" when x"87",
		x"0B" when x"88",
		x"09" when x"89",
		x"0F" when x"8A",
		x"0D" when x"8B",
		x"03" when x"8C",
		x"01" when x"8D",
		x"07" when x"8E",
		x"05" when x"8F",
		x"3B" when x"90",
		x"39" when x"91",
		x"3F" when x"92",
		x"3D" when x"93",
		x"33" when x"94",
		x"31" when x"95",
		x"37" when x"96",
		x"35" when x"97",
		x"2B" when x"98",
		x"29" when x"99",
		x"2F" when x"9A",
		x"2D" when x"9B",
		x"23" when x"9C",
		x"21" when x"9D",
		x"27" when x"9E",
		x"25" when x"9F",
		x"5B" when x"A0",
		x"59" when x"A1",
		x"5F" when x"A2",
		x"5D" when x"A3",
		x"53" when x"A4",
		x"51" when x"A5",
		x"57" when x"A6",
		x"55" when x"A7",
		x"4B" when x"A8",
		x"49" when x"A9",
		x"4F" when x"AA",
		x"4D" when x"AB",
		x"43" when x"AC",
		x"41" when x"AD",
		x"47" when x"AE",
		x"45" when x"AF",
		x"7B" when x"B0",
		x"79" when x"B1",
		x"7F" when x"B2",
		x"7D" when x"B3",
		x"73" when x"B4",
		x"71" when x"B5",
		x"77" when x"B6",
		x"75" when x"B7",
		x"6B" when x"B8",
		x"69" when x"B9",
		x"6F" when x"BA",
		x"6D" when x"BB",
		x"63" when x"BC",
		x"61" when x"BD",
		x"67" when x"BE",
		x"65" when x"BF",
		x"9B" when x"C0",
		x"99" when x"C1",
		x"9F" when x"C2",
		x"9D" when x"C3",
		x"93" when x"C4",
		x"91" when x"C5",
		x"97" when x"C6",
		x"95" when x"C7",
		x"8B" when x"C8",
		x"89" when x"C9",
		x"8F" when x"CA",
		x"8D" when x"CB",
		x"83" when x"CC",
		x"81" when x"CD",
		x"87" when x"CE",
		x"85" when x"CF",
		x"BB" when x"D0",
		x"B9" when x"D1",
		x"BF" when x"D2",
		x"BD" when x"D3",
		x"B3" when x"D4",
		x"B1" when x"D5",
		x"B7" when x"D6",
		x"B5" when x"D7",
		x"AB" when x"D8",
		x"A9" when x"D9",
		x"AF" when x"DA",
		x"AD" when x"DB",
		x"A3" when x"DC",
		x"A1" when x"DD",
		x"A7" when x"DE",
		x"A5" when x"DF",
		x"DB" when x"E0",
		x"D9" when x"E1",
		x"DF" when x"E2",
		x"DD" when x"E3",
		x"D3" when x"E4",
		x"D1" when x"E5",
		x"D7" when x"E6",
		x"D5" when x"E7",
		x"CB" when x"E8",
		x"C9" when x"E9",
		x"CF" when x"EA",
		x"CD" when x"EB",
		x"C3" when x"EC",
		x"C1" when x"ED",
		x"C7" when x"EE",
		x"C5" when x"EF",
		x"FB" when x"F0",
		x"F9" when x"F1",
		x"FF" when x"F2",
		x"FD" when x"F3",
		x"F3" when x"F4",
		x"F1" when x"F5",
		x"F7" when x"F6",
		x"F5" when x"F7",
		x"EB" when x"F8",
		x"E9" when x"F9",
		x"EF" when x"FA",
		x"ED" when x"FB",
		x"E3" when x"FC",
		x"E1" when x"FD",
		x"E7" when x"FE",
		x"E5" when x"FF",
		x"00" when others;

end Behavioral;

